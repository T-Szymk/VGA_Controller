/*******************************************************************************
-- Title      : VGA Line Buffer Controller
-- Project    : VGA Controller
********************************************************************************
-- File       : line_buff_ctrl.sv
-- Author(s)  : Thomas Szymkowiak
-- Company    : TUNI
-- Created    : 2022-08-21
-- Design     : line_buff_ctrl
-- Platform   : -
-- Standard   : SystemVerilog '17
********************************************************************************
-- Description: VGA line buffer controller model written in SV
********************************************************************************
-- Revisions:
-- Date        Version  Author  Description
-- 2022-08-21  1.0      TZS     Created
*******************************************************************************/